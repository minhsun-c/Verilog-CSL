`include "src/CLA.v"

module tb;
    reg [3:0] A, B;
    wire [3:0] Sum;
    wire Cout;

    CLA_Adder4 CA(
        .Cout(Cout),
        .Sum(Sum),
        .A(A), 
        .B(B),
        .Cin(1'b0)
    );

    initial begin
        $monitor(
            "[%03g] %04b + %04b = %b%04b",
            $time, A, B, Cout, Sum
        );
        // for (integer i=0; i<16; i=i+1) begin
        //     for (integer j=0; j<16; j=j+1) begin
        //         #1 A = i; B = j; 
        //         $display(
        //             "[%3g] %04b + %04b = %b%04b",
        //             $time, A, B, Cout, Sum
        //         );
        //     end
        // end
        #1 A = 4'd0; B = 4'd0;
		#1 A = 4'd0; B = 4'd1;
		#1 A = 4'd0; B = 4'd2;
		#1 A = 4'd0; B = 4'd3;
		#1 A = 4'd0; B = 4'd4;
		#1 A = 4'd0; B = 4'd5;
		#1 A = 4'd0; B = 4'd6;
		#1 A = 4'd0; B = 4'd7;
		#1 A = 4'd0; B = 4'd8;
		#1 A = 4'd0; B = 4'd9;
		#1 A = 4'd0; B = 4'd10;
		#1 A = 4'd0; B = 4'd11;
		#1 A = 4'd0; B = 4'd12;
		#1 A = 4'd0; B = 4'd13;
		#1 A = 4'd0; B = 4'd14;
		#1 A = 4'd0; B = 4'd15;
		#1 A = 4'd1; B = 4'd0;
		#1 A = 4'd1; B = 4'd1;
		#1 A = 4'd1; B = 4'd2;
		#1 A = 4'd1; B = 4'd3;
		#1 A = 4'd1; B = 4'd4;
		#1 A = 4'd1; B = 4'd5;
		#1 A = 4'd1; B = 4'd6;
		#1 A = 4'd1; B = 4'd7;
		#1 A = 4'd1; B = 4'd8;
		#1 A = 4'd1; B = 4'd9;
		#1 A = 4'd1; B = 4'd10;
		#1 A = 4'd1; B = 4'd11;
		#1 A = 4'd1; B = 4'd12;
		#1 A = 4'd1; B = 4'd13;
		#1 A = 4'd1; B = 4'd14;
		#1 A = 4'd1; B = 4'd15;
		#1 A = 4'd2; B = 4'd0;
		#1 A = 4'd2; B = 4'd1;
		#1 A = 4'd2; B = 4'd2;
		#1 A = 4'd2; B = 4'd3;
		#1 A = 4'd2; B = 4'd4;
		#1 A = 4'd2; B = 4'd5;
		#1 A = 4'd2; B = 4'd6;
		#1 A = 4'd2; B = 4'd7;
		#1 A = 4'd2; B = 4'd8;
		#1 A = 4'd2; B = 4'd9;
		#1 A = 4'd2; B = 4'd10;
		#1 A = 4'd2; B = 4'd11;
		#1 A = 4'd2; B = 4'd12;
		#1 A = 4'd2; B = 4'd13;
		#1 A = 4'd2; B = 4'd14;
		#1 A = 4'd2; B = 4'd15;
		#1 A = 4'd3; B = 4'd0;
		#1 A = 4'd3; B = 4'd1;
		#1 A = 4'd3; B = 4'd2;
		#1 A = 4'd3; B = 4'd3;
		#1 A = 4'd3; B = 4'd4;
		#1 A = 4'd3; B = 4'd5;
		#1 A = 4'd3; B = 4'd6;
		#1 A = 4'd3; B = 4'd7;
		#1 A = 4'd3; B = 4'd8;
		#1 A = 4'd3; B = 4'd9;
		#1 A = 4'd3; B = 4'd10;
		#1 A = 4'd3; B = 4'd11;
		#1 A = 4'd3; B = 4'd12;
		#1 A = 4'd3; B = 4'd13;
		#1 A = 4'd3; B = 4'd14;
		#1 A = 4'd3; B = 4'd15;
		#1 A = 4'd4; B = 4'd0;
		#1 A = 4'd4; B = 4'd1;
		#1 A = 4'd4; B = 4'd2;
		#1 A = 4'd4; B = 4'd3;
		#1 A = 4'd4; B = 4'd4;
		#1 A = 4'd4; B = 4'd5;
		#1 A = 4'd4; B = 4'd6;
		#1 A = 4'd4; B = 4'd7;
		#1 A = 4'd4; B = 4'd8;
		#1 A = 4'd4; B = 4'd9;
		#1 A = 4'd4; B = 4'd10;
		#1 A = 4'd4; B = 4'd11;
		#1 A = 4'd4; B = 4'd12;
		#1 A = 4'd4; B = 4'd13;
		#1 A = 4'd4; B = 4'd14;
		#1 A = 4'd4; B = 4'd15;
		#1 A = 4'd5; B = 4'd0;
		#1 A = 4'd5; B = 4'd1;
		#1 A = 4'd5; B = 4'd2;
		#1 A = 4'd5; B = 4'd3;
		#1 A = 4'd5; B = 4'd4;
		#1 A = 4'd5; B = 4'd5;
		#1 A = 4'd5; B = 4'd6;
		#1 A = 4'd5; B = 4'd7;
		#1 A = 4'd5; B = 4'd8;
		#1 A = 4'd5; B = 4'd9;
		#1 A = 4'd5; B = 4'd10;
		#1 A = 4'd5; B = 4'd11;
		#1 A = 4'd5; B = 4'd12;
		#1 A = 4'd5; B = 4'd13;
		#1 A = 4'd5; B = 4'd14;
		#1 A = 4'd5; B = 4'd15;
		#1 A = 4'd6; B = 4'd0;
		#1 A = 4'd6; B = 4'd1;
		#1 A = 4'd6; B = 4'd2;
		#1 A = 4'd6; B = 4'd3;
		#1 A = 4'd6; B = 4'd4;
		#1 A = 4'd6; B = 4'd5;
		#1 A = 4'd6; B = 4'd6;
		#1 A = 4'd6; B = 4'd7;
		#1 A = 4'd6; B = 4'd8;
		#1 A = 4'd6; B = 4'd9;
		#1 A = 4'd6; B = 4'd10;
		#1 A = 4'd6; B = 4'd11;
		#1 A = 4'd6; B = 4'd12;
		#1 A = 4'd6; B = 4'd13;
		#1 A = 4'd6; B = 4'd14;
		#1 A = 4'd6; B = 4'd15;
		#1 A = 4'd7; B = 4'd0;
		#1 A = 4'd7; B = 4'd1;
		#1 A = 4'd7; B = 4'd2;
		#1 A = 4'd7; B = 4'd3;
		#1 A = 4'd7; B = 4'd4;
		#1 A = 4'd7; B = 4'd5;
		#1 A = 4'd7; B = 4'd6;
		#1 A = 4'd7; B = 4'd7;
		#1 A = 4'd7; B = 4'd8;
		#1 A = 4'd7; B = 4'd9;
		#1 A = 4'd7; B = 4'd10;
		#1 A = 4'd7; B = 4'd11;
		#1 A = 4'd7; B = 4'd12;
		#1 A = 4'd7; B = 4'd13;
		#1 A = 4'd7; B = 4'd14;
		#1 A = 4'd7; B = 4'd15;
		#1 A = 4'd8; B = 4'd0;
		#1 A = 4'd8; B = 4'd1;
		#1 A = 4'd8; B = 4'd2;
		#1 A = 4'd8; B = 4'd3;
		#1 A = 4'd8; B = 4'd4;
		#1 A = 4'd8; B = 4'd5;
		#1 A = 4'd8; B = 4'd6;
		#1 A = 4'd8; B = 4'd7;
		#1 A = 4'd8; B = 4'd8;
		#1 A = 4'd8; B = 4'd9;
		#1 A = 4'd8; B = 4'd10;
		#1 A = 4'd8; B = 4'd11;
		#1 A = 4'd8; B = 4'd12;
		#1 A = 4'd8; B = 4'd13;
		#1 A = 4'd8; B = 4'd14;
		#1 A = 4'd8; B = 4'd15;
		#1 A = 4'd9; B = 4'd0;
		#1 A = 4'd9; B = 4'd1;
		#1 A = 4'd9; B = 4'd2;
		#1 A = 4'd9; B = 4'd3;
		#1 A = 4'd9; B = 4'd4;
		#1 A = 4'd9; B = 4'd5;
		#1 A = 4'd9; B = 4'd6;
		#1 A = 4'd9; B = 4'd7;
		#1 A = 4'd9; B = 4'd8;
		#1 A = 4'd9; B = 4'd9;
		#1 A = 4'd9; B = 4'd10;
		#1 A = 4'd9; B = 4'd11;
		#1 A = 4'd9; B = 4'd12;
		#1 A = 4'd9; B = 4'd13;
		#1 A = 4'd9; B = 4'd14;
		#1 A = 4'd9; B = 4'd15;
		#1 A = 4'd10; B = 4'd0;
		#1 A = 4'd10; B = 4'd1;
		#1 A = 4'd10; B = 4'd2;
		#1 A = 4'd10; B = 4'd3;
		#1 A = 4'd10; B = 4'd4;
		#1 A = 4'd10; B = 4'd5;
		#1 A = 4'd10; B = 4'd6;
		#1 A = 4'd10; B = 4'd7;
		#1 A = 4'd10; B = 4'd8;
		#1 A = 4'd10; B = 4'd9;
		#1 A = 4'd10; B = 4'd10;
		#1 A = 4'd10; B = 4'd11;
		#1 A = 4'd10; B = 4'd12;
		#1 A = 4'd10; B = 4'd13;
		#1 A = 4'd10; B = 4'd14;
		#1 A = 4'd10; B = 4'd15;
		#1 A = 4'd11; B = 4'd0;
		#1 A = 4'd11; B = 4'd1;
		#1 A = 4'd11; B = 4'd2;
		#1 A = 4'd11; B = 4'd3;
		#1 A = 4'd11; B = 4'd4;
		#1 A = 4'd11; B = 4'd5;
		#1 A = 4'd11; B = 4'd6;
		#1 A = 4'd11; B = 4'd7;
		#1 A = 4'd11; B = 4'd8;
		#1 A = 4'd11; B = 4'd9;
		#1 A = 4'd11; B = 4'd10;
		#1 A = 4'd11; B = 4'd11;
		#1 A = 4'd11; B = 4'd12;
		#1 A = 4'd11; B = 4'd13;
		#1 A = 4'd11; B = 4'd14;
		#1 A = 4'd11; B = 4'd15;
		#1 A = 4'd12; B = 4'd0;
		#1 A = 4'd12; B = 4'd1;
		#1 A = 4'd12; B = 4'd2;
		#1 A = 4'd12; B = 4'd3;
		#1 A = 4'd12; B = 4'd4;
		#1 A = 4'd12; B = 4'd5;
		#1 A = 4'd12; B = 4'd6;
		#1 A = 4'd12; B = 4'd7;
		#1 A = 4'd12; B = 4'd8;
		#1 A = 4'd12; B = 4'd9;
		#1 A = 4'd12; B = 4'd10;
		#1 A = 4'd12; B = 4'd11;
		#1 A = 4'd12; B = 4'd12;
		#1 A = 4'd12; B = 4'd13;
		#1 A = 4'd12; B = 4'd14;
		#1 A = 4'd12; B = 4'd15;
		#1 A = 4'd13; B = 4'd0;
		#1 A = 4'd13; B = 4'd1;
		#1 A = 4'd13; B = 4'd2;
		#1 A = 4'd13; B = 4'd3;
		#1 A = 4'd13; B = 4'd4;
		#1 A = 4'd13; B = 4'd5;
		#1 A = 4'd13; B = 4'd6;
		#1 A = 4'd13; B = 4'd7;
		#1 A = 4'd13; B = 4'd8;
		#1 A = 4'd13; B = 4'd9;
		#1 A = 4'd13; B = 4'd10;
		#1 A = 4'd13; B = 4'd11;
		#1 A = 4'd13; B = 4'd12;
		#1 A = 4'd13; B = 4'd13;
		#1 A = 4'd13; B = 4'd14;
		#1 A = 4'd13; B = 4'd15;
		#1 A = 4'd14; B = 4'd0;
		#1 A = 4'd14; B = 4'd1;
		#1 A = 4'd14; B = 4'd2;
		#1 A = 4'd14; B = 4'd3;
		#1 A = 4'd14; B = 4'd4;
		#1 A = 4'd14; B = 4'd5;
		#1 A = 4'd14; B = 4'd6;
		#1 A = 4'd14; B = 4'd7;
		#1 A = 4'd14; B = 4'd8;
		#1 A = 4'd14; B = 4'd9;
		#1 A = 4'd14; B = 4'd10;
		#1 A = 4'd14; B = 4'd11;
		#1 A = 4'd14; B = 4'd12;
		#1 A = 4'd14; B = 4'd13;
		#1 A = 4'd14; B = 4'd14;
		#1 A = 4'd14; B = 4'd15;
		#1 A = 4'd15; B = 4'd0;
		#1 A = 4'd15; B = 4'd1;
		#1 A = 4'd15; B = 4'd2;
		#1 A = 4'd15; B = 4'd3;
		#1 A = 4'd15; B = 4'd4;
		#1 A = 4'd15; B = 4'd5;
		#1 A = 4'd15; B = 4'd6;
		#1 A = 4'd15; B = 4'd7;
		#1 A = 4'd15; B = 4'd8;
		#1 A = 4'd15; B = 4'd9;
		#1 A = 4'd15; B = 4'd10;
		#1 A = 4'd15; B = 4'd11;
		#1 A = 4'd15; B = 4'd12;
		#1 A = 4'd15; B = 4'd13;
		#1 A = 4'd15; B = 4'd14;
		#1 A = 4'd15; B = 4'd15;

        

    end
endmodule