`ifndef _FINITE_STATE_MACHINE 
`define _FINITE_STATE_MACHINE

/*
    state: 
*/
module FSM (
    output reg out,
    input areset,
    input [1:0] data, // data for reseting the fsm
    input in
);
    always @() begin
        
    end
    
endmodule

`endif 